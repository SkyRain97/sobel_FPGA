`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2021/07/12 17:25:15
// Design Name: 
// Module Name: sobel_data_buffer_mod_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

`define clk_period 10

module sobel_data_buffer_mod_tb();
reg         clk, rst, done_i;
reg  [7:0]  grayscale_i;
wire [7:0]  d0_o, d1_o, d2_o, d3_o, d4_o, d5_o, d6_o, d7_o, d8_o;
wire        done_o;

sobel_data_buffer_mod #(.ROWS(5), .COLS(6)) SOBEL_DATA_BUFFER_MOD(
    .clk(clk),
    .rst(rst),
    .done_i(done_i),
    .grayscale_i(grayscale_i),

    .d0_o(d0_o), .d1_o(d1_o), .d2_o(d2_o), .d3_o(d3_o), .d4_o(d4_o), .d5_o(d5_o), .d6_o(d6_o), .d7_o(d7_o), .d8_o(d8_o),
    .done_o(done_o)
);

initial clk = 1'b1;
always #(`clk_period/2) clk = ~clk;

integer i;

initial begin
    rst = 1'b1;
    grayscale_i = 8'b0;
    done_i = 1'b0;

    #(`clk_period);
    rst = 1'b0;
    done_i = 1'b1;

    for(i = 1; i < 36; i = i + 1) begin
        grayscale_i = i;
        #(`clk_period);
    end

    done_i = 1'b0;

    #(`clk_period);
    $stop;



end
endmodule
